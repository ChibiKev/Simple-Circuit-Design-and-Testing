library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_8To3Encoder is
    port(
        Chen_Kevin_O1   : out    vl_logic;
        Chen_Kevin_I8   : in     vl_logic;
        Chen_Kevin_I4   : in     vl_logic;
        Chen_Kevin_I2   : in     vl_logic;
        Chen_Kevin_I6   : in     vl_logic;
        Chen_Kevin_O2   : out    vl_logic;
        Chen_Kevin_I3   : in     vl_logic;
        Chen_Kevin_I7   : in     vl_logic;
        Chen_Kevin_O3   : out    vl_logic;
        Chen_Kevin_I5   : in     vl_logic;
        Chen_Kevin_I1   : in     vl_logic
    );
end Chen_Kevin_8To3Encoder;
