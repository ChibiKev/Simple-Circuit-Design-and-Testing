library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_8T3Encoder_vlg_sample_tst is
    port(
        Chen_Kevin_I1   : in     vl_logic;
        Chen_Kevin_I2   : in     vl_logic;
        Chen_Kevin_I3   : in     vl_logic;
        Chen_Kevin_I4   : in     vl_logic;
        Chen_Kevin_I5   : in     vl_logic;
        Chen_Kevin_I6   : in     vl_logic;
        Chen_Kevin_I7   : in     vl_logic;
        Chen_Kevin_I8   : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Chen_Kevin_8T3Encoder_vlg_sample_tst;
