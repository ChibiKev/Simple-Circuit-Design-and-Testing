library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_8T3Encoder_vlg_check_tst is
    port(
        Chen_Kevin_O1   : in     vl_logic;
        Chen_Kevin_O2   : in     vl_logic;
        Chen_Kevin_O3   : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_8T3Encoder_vlg_check_tst;
