library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_1BitFullAdderUsing1BitHalfAdderAsAComponent_vlg_sample_tst is
    port(
        Chen_Kevin_Cin  : in     vl_logic;
        Chen_Kevin_I1   : in     vl_logic;
        Chen_Kevin_I2   : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Chen_Kevin_1BitFullAdderUsing1BitHalfAdderAsAComponent_vlg_sample_tst;
