library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_1BitFullAdderUsing1BitHalfAdderAsAComponent_vlg_check_tst is
    port(
        Chen_Kevin_Cout : in     vl_logic;
        Chen_Kevin_S    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_1BitFullAdderUsing1BitHalfAdderAsAComponent_vlg_check_tst;
