library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_SimpleCircuit_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_SimpleCircuit_vlg_check_tst;
