library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_3T8Decoder is
    port(
        Chen_Kevin_I1   : in     vl_logic;
        Chen_Kevin_I2   : in     vl_logic;
        Chen_Kevin_I3   : in     vl_logic;
        Chen_Kevin_O1   : out    vl_logic;
        Chen_Kevin_O2   : out    vl_logic;
        Chen_Kevin_O3   : out    vl_logic;
        Chen_Kevin_O4   : out    vl_logic;
        Chen_Kevin_O5   : out    vl_logic;
        Chen_Kevin_O6   : out    vl_logic;
        Chen_Kevin_O7   : out    vl_logic;
        Chen_Kevin_O8   : out    vl_logic
    );
end Chen_Kevin_3T8Decoder;
