library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Mux2to1_vlg_vec_tst is
end Chen_Kevin_Mux2to1_vlg_vec_tst;
