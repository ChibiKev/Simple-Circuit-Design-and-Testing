library verilog;
use verilog.vl_types.all;
entity DecoderLPM_vlg_vec_tst is
end DecoderLPM_vlg_vec_tst;
