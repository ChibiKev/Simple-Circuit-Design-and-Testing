library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_FullAdderLPM_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        result          : in     vl_logic_vector(0 downto 0);
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_FullAdderLPM_vlg_check_tst;
