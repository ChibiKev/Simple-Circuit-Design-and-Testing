library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Mux2to1 is
    port(
        Chen_Kevin_M    : out    vl_logic;
        Chen_Kevin_S    : in     vl_logic;
        Chen_Kevin_Y    : in     vl_logic;
        Chen_Kevin_X    : in     vl_logic
    );
end Chen_Kevin_Mux2to1;
