library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Mux2to1_vlg_check_tst is
    port(
        Chen_Kevin_M    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_Mux2to1_vlg_check_tst;
