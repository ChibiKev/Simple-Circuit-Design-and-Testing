library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_SimpleCircuit is
    port(
        f               : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end Chen_Kevin_SimpleCircuit;
