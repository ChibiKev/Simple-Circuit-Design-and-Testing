library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_Mux2to1_vlg_sample_tst is
    port(
        Chen_Kevin_S    : in     vl_logic;
        Chen_Kevin_X    : in     vl_logic;
        Chen_Kevin_Y    : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Chen_Kevin_Mux2to1_vlg_sample_tst;
