library verilog;
use verilog.vl_types.all;
entity DecoderLPM_vlg_check_tst is
    port(
        eq0             : in     vl_logic;
        eq1             : in     vl_logic;
        eq2             : in     vl_logic;
        eq3             : in     vl_logic;
        eq4             : in     vl_logic;
        eq5             : in     vl_logic;
        eq6             : in     vl_logic;
        eq7             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DecoderLPM_vlg_check_tst;
