library verilog;
use verilog.vl_types.all;
entity Chen_Kevin_MuxLPM_vlg_check_tst is
    port(
        result          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Chen_Kevin_MuxLPM_vlg_check_tst;
